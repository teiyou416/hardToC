module out;
initial begin $display("Hello"); $finish;end
endmodule
